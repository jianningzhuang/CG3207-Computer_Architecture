
----------------------------------------------------------------
-- Instruction Memory
----------------------------------------------------------------
constant INSTR_MEM : MEM_128x32 := (		x"159F11F8", 
											x"359F21F8", 
											x"559F31F8", 
											x"759F4204", 
											x"E59F5214", 
											x"E59F6200", 
											x"E59F720C", 
											x"E59F8208", 
											x"E59FB1FC", 
											x"E38CC0FF", 
											x"E59FD1F8", 
											x"E09DC0AC", 
											x"600CC006", 
											x"415C000C", 
											x"017D008D", 
											x"2591C004", 
											x"2502C004", 
											x"225BB001", 
											x"CAFFFFF5", 
											x"EAFFFFFF", 
											x"E35500FA", 
											x"D59F61D4", 
											x"E35500E1", 
											x"C5846000", 
											x"E35500E1", 
											x"D59F61C8", 
											x"E35500C8", 
											x"C5846000", 
											x"E35500C8", 
											x"D59F61BC", 
											x"E35500AF", 
											x"C5846000", 
											x"E35500AF", 
											x"D59F6190", 
											x"D5846000", 
											x"E5936000", 
											x"E58F5768", 
											x"E3560004", 
											x"059F7760", 
											x"E3560001", 
											x"059F8758", 
											x"E3560005", 
											x"059F7750", 
											x"059F874C", 
											x"E2555001", 
											x"1AFFFFE5", 
											x"EAFFFFFF", 
											x"E5936000", 
											x"E58F5738", 
											x"E3560004", 
											x"059F7730", 
											x"E3560001", 
											x"059F8728", 
											x"E3560005", 
											x"059F7720", 
											x"059F871C", 
											x"E2855001", 
											x"E3550064", 
											x"1AFFFFF3", 
											x"EAFFFFFF", 
											x"E1570008", 
											x"C59F6144", 
											x"C5846000", 
											x"B59F6138", 
											x"B5846000", 
											x"059F6138", 
											x"05846000", 
											x"EAFFFFFF", 
											x"E5926000", 
											x"E5816000", 
											x"EAFFFFFC", 
											x"EAFFFFFE", 
											others => x"00000000");

----------------------------------------------------------------
-- Data (Constant) Memory
----------------------------------------------------------------
constant DATA_CONST_MEM : MEM_128x32 := (	x"00000C00", 
											x"00000C04", 
											x"00000C08", 
											x"00000C0C", 
											x"00000C10", 
											x"00000C14", 
											x"00000C18", 
											x"00000000", 
											x"000000FF", 
											x"00000064", 
											x"7FFFFFFF", 
											x"000000FA", 
											x"01000100", 
											x"00900090", 
											x"00800080", 
											x"AAAAAAAA", 
											x"BBBBBBBB", 
											x"AAAABBBB", 
											x"00000800", 
											x"ABCD1234", 
											x"65570A0D", 
											x"6D6F636C", 
											x"6F742065", 
											x"33474320", 
											x"2E373032", 
											x"000A0D2E", 
											x"00000250", 
											others => x"00000000");

